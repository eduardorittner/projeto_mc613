module cobra (
  input clk,
  input up,
  input down,
  input left,
  input right,
  output next_pos
);

endmodule
